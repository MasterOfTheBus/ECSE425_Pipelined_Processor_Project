LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY ALUController IS
	PORT(	
		opcode		: IN std_logic_vector(5 DOWNTO 0);
		
		-- EX Stage
		RegDst		: OUT std_logic;
		ALUOp		: OUT std_logic_vector(1 DOWNTO 0);
		ALUSrc		: OUT std_logic;
		-- MEM Stage
		Branch		: OUT std_logic;
		MemRead		: OUT std_logic;
		MemWrite	: OUT std_logic;
		-- WB Stage
		RegWrite	: OUT std_logic;
		MemtoReg	: OUT std_logic
	);
	END ENTITY;
	
ARCHITECTURE behavior OF ALUController IS
	SIGNAL ctrl_matrix: std_logic_vector(8 downto 0);
BEGIN
	PROCESS(opcode) 
		BEGIN
		CASE opcode IS
			WHEN "000000" => ctrl_matrix <= "100100010"; -- R-type
            WHEN "100011" => ctrl_matrix <= "011110000"; -- lw
            WHEN "101011" => ctrl_matrix <= "010001000"; -- sw
            WHEN "000100" => ctrl_matrix <= "000000101"; -- beq
            
			-- WHEN "001000" => ctrl_matrix <= "011000000"; -- addi
            -- WHEN "000010" => ctrl_matrix <= "000000100"; -- j
            -- WHEN "000011" => ctrl_matrix <= "001000001"; -- jal
            -- WHEN "001001" => ctrl_matrix <= "011000001"; -- subi
            WHEN OTHERS   => ctrl_matrix <= "---------";
		END CASE;
		
	RegDst		<= ctrl_matrix(8);
	ALUSrc		<= ctrl_matrix(7);
	MemtoReg	<= ctrl_matrix(6);
	RegWrite	<= ctrl_matrix(5);
	MemWrite	<= ctrl_matrix(4);
	MemRead		<= ctrl_matrix(3);
	Branch		<= ctrl_matrix(2);
	ALUOp		<= ctrl_matrix(1 DOWNTO 0);
	END PROCESS;	
END behavior;